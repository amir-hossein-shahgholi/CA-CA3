module shl2_32b(input [31:0] IN,output [31:0] out);
    assign out = IN << 2;
endmodule